magic
tech sky130A
magscale 1 2
timestamp 1762969946
<< error_s >>
rect 1605 1417 1663 1423
rect 1605 1383 1617 1417
rect 1605 1377 1663 1383
rect 1036 809 1071 843
rect 1459 826 1493 844
rect 1037 790 1071 809
rect 867 741 925 747
rect 298 697 333 731
rect 721 714 755 732
rect 299 678 333 697
rect 129 629 187 635
rect 129 595 141 629
rect 129 589 187 595
rect 129 119 187 125
rect 129 85 141 119
rect 129 79 187 85
rect 318 -17 333 678
rect 352 644 387 678
rect 352 -17 386 644
rect 498 576 556 582
rect 498 542 510 576
rect 498 536 556 542
rect 498 66 556 72
rect 498 32 510 66
rect 498 26 556 32
rect 352 -51 367 -17
rect 685 -70 755 714
rect 867 707 879 741
rect 867 701 925 707
rect 867 13 925 19
rect 867 -21 879 13
rect 867 -27 925 -21
rect 685 -106 738 -70
rect 1056 -123 1071 790
rect 1090 756 1125 790
rect 1090 -123 1124 756
rect 1236 688 1294 694
rect 1236 654 1248 688
rect 1236 648 1294 654
rect 1236 -40 1294 -34
rect 1236 -74 1248 -40
rect 1236 -80 1294 -74
rect 1090 -157 1105 -123
rect 1423 -176 1493 826
rect 1605 -93 1663 -87
rect 1605 -127 1617 -93
rect 1605 -133 1663 -127
rect 1423 -212 1476 -176
use sky130_fd_pr__nfet_01v8_ATLS57  XM1
timestamp 1762969946
transform 1 0 158 0 1 357
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_XGSNAL  XM2
timestamp 1762969946
transform 1 0 896 0 1 360
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_ATLS57  XM3
timestamp 1762969946
transform 1 0 527 0 1 304
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_XGSNAL  XM4
timestamp 1762969946
transform 1 0 1265 0 1 307
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_KBNS5F  XM5
timestamp 1762969946
transform 1 0 1634 0 1 645
box -211 -910 211 910
<< end >>
