magic
tech sky130A
magscale 1 2
timestamp 1764122104
<< error_p >>
rect -29 572 29 578
rect -29 538 -17 572
rect -29 532 29 538
rect -29 -538 29 -532
rect -29 -572 -17 -538
rect -29 -578 29 -572
<< pwell >>
rect -211 -710 211 710
<< nmos >>
rect -15 -500 15 500
<< ndiff >>
rect -73 488 -15 500
rect -73 -488 -61 488
rect -27 -488 -15 488
rect -73 -500 -15 -488
rect 15 488 73 500
rect 15 -488 27 488
rect 61 -488 73 488
rect 15 -500 73 -488
<< ndiffc >>
rect -61 -488 -27 488
rect 27 -488 61 488
<< psubdiff >>
rect -175 640 -79 674
rect 79 640 175 674
rect -175 578 -141 640
rect 141 578 175 640
rect -175 -640 -141 -578
rect 141 -640 175 -578
rect -175 -674 -79 -640
rect 79 -674 175 -640
<< psubdiffcont >>
rect -79 640 79 674
rect -175 -578 -141 578
rect 141 -578 175 578
rect -79 -674 79 -640
<< poly >>
rect -33 572 33 588
rect -33 538 -17 572
rect 17 538 33 572
rect -33 522 33 538
rect -15 500 15 522
rect -15 -522 15 -500
rect -33 -538 33 -522
rect -33 -572 -17 -538
rect 17 -572 33 -538
rect -33 -588 33 -572
<< polycont >>
rect -17 538 17 572
rect -17 -572 17 -538
<< locali >>
rect -175 640 -79 674
rect 79 640 175 674
rect -175 578 -141 640
rect 141 578 175 640
rect -33 538 -17 572
rect 17 538 33 572
rect -61 488 -27 504
rect -61 -504 -27 -488
rect 27 488 61 504
rect 27 -504 61 -488
rect -33 -572 -17 -538
rect 17 -572 33 -538
rect -175 -640 -141 -578
rect 141 -640 175 -578
rect -175 -674 -79 -640
rect 79 -674 175 -640
<< viali >>
rect -17 538 17 572
rect -61 -488 -27 488
rect 27 -488 61 488
rect -17 -572 17 -538
<< metal1 >>
rect -29 572 29 578
rect -29 538 -17 572
rect 17 538 29 572
rect -29 532 29 538
rect -67 488 -21 500
rect -67 -488 -61 488
rect -27 -488 -21 488
rect -67 -500 -21 -488
rect 21 488 67 500
rect 21 -488 27 488
rect 61 -488 67 488
rect 21 -500 67 -488
rect -29 -538 29 -532
rect -29 -572 -17 -538
rect 17 -572 29 -538
rect -29 -578 29 -572
<< properties >>
string FIXED_BBOX -158 -657 158 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
