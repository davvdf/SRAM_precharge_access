magic
tech sky130A
magscale 1 2
timestamp 1764873183
<< locali >>
rect 299 85 437 119
rect 719 85 857 119
<< metal1 >>
rect 141 2195 1015 2230
rect 141 1195 175 2195
rect 981 1194 1015 2195
rect 185 759 551 959
rect 605 760 971 960
rect 40 380 141 399
rect 40 319 80 380
rect 140 319 141 380
rect 40 299 141 319
rect 1013 381 1114 400
rect 1073 320 1114 381
rect 1013 300 1114 320
rect 141 85 1015 119
<< via1 >>
rect 80 319 140 380
rect 1013 320 1073 381
<< metal2 >>
rect 40 381 1114 399
rect 40 380 1013 381
rect 40 319 80 380
rect 140 320 1013 380
rect 1073 320 1114 381
rect 140 319 1114 320
rect 40 300 1114 319
use sky130_fd_pr__nfet_01v8_66AFG5  sky130_fd_pr__nfet_01v8_66AFG5_0
timestamp 1764122104
transform 1 0 578 0 1 1157
box -211 -1210 211 1210
use sky130_fd_pr__nfet_01v8_GV8PYF  sky130_fd_pr__nfet_01v8_GV8PYF_0
timestamp 1764122104
transform 1 0 158 0 1 657
box -211 -710 211 710
use sky130_fd_pr__nfet_01v8_GV8PYF  sky130_fd_pr__nfet_01v8_GV8PYF_1
timestamp 1764122104
transform 1 0 998 0 1 657
box -211 -710 211 710
<< labels >>
flabel metal1 185 759 551 959 0 FreeSans 160 0 0 0 BL
port 2 nsew
flabel space 599 760 977 960 0 FreeSans 160 0 0 0 BL_N
port 3 nsew
flabel metal1 141 2195 1015 2230 0 FreeSans 160 0 0 0 CLK
port 1 nsew
flabel metal1 141 85 1015 119 0 FreeSans 160 0 0 0 VSS
port 5 nsew
flabel metal2 40 300 1114 399 0 FreeSans 160 0 0 0 0.5VDD
port 6 nsew
<< end >>
