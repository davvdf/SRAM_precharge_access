** sch_path: /home/david/Documents/SRAM_precharge_access/analog/schematics/trans_gate_tb.sch
**.subckt trans_gate_tb
V3 clk GND PULSE(0 1.8 0n 0.2n 0.2n 7.5n 15.15n)
x2 clk VGND VNB VPB VPWR net3 sky130_fd_sc_hd__clkinv_1
V4 net1 GND DC 0.9 AC 0.001
CBLB BL_N GND 300f m=1
CBL BL GND 300f m=1
x1 net3 BL_N BL net2 net1 clk precharge_trans_gate
V1 net2 GND DC 1.8 AC 0.001
**** begin user architecture code

.include "/home/david/.volare/volare/sky130/versions/fa87f8f4bbcc7255b6f0c0fb506960f531ae2392/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice"

.ic V(BL)=0.895 V(BL_n)=0.905V
.control
* Nested loops for all corners
foreach temp_val -40 27 125
  foreach vdd_val 1.79 1.8 1.81
      reset
      alter V1 = $vdd_val
      set temp = $temp_val


      tran 0.001n 0.5n
      let new_val=abs(V(BL_n)-V(BL))
      meas tran t_pch WHEN new_val=0.002 CROSS=1

      echo "T=$temp_val, VDD=$vdd_val, t_pch=$&t_pch"
    * >> smallest_diff.txt
    end
  end
end
plot tran1.new_val tran2.new_val tran3.new_val tran4.new_val tran5.new_val tran6.new_val
+ tran7.new_val tran8.new_val tran9.new_val
rusage all
.endc
.noise v(BL) V4 dec 10 1 66MEG


.param mc_mm_switch=1
.param mc_pr_switch=0
.include /home/david/.volare/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/david/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/david/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/david/.volare/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  precharge_trans_gate.sym # of pins=6
** sym_path: /home/david/Documents/SRAM_precharge_access/analog/schematics/precharge_trans_gate.sym
** sch_path: /home/david/Documents/SRAM_precharge_access/analog/schematics/precharge_trans_gate.sch
.subckt precharge_trans_gate clk_n BL_N BL VDD VDD_div2 clk
*.ipin VDD_div2
*.ipin clk_n
*.ipin clk
*.iopin BL
*.iopin BL_N
*.ipin VDD
XM1 VDD_div2 clk BL GND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 BL_N clk VDD_div2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 VDD_div2 clk_n BL VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 BL_N clk_n VDD_div2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 BL clk BL_N GND sky130_fd_pr__nfet_01v8 L=0.15 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
