magic
tech sky130A
magscale 1 2
timestamp 1763573990
<< error_s >>
rect 1422 2584 1480 2590
rect 1422 2550 1434 2584
rect 1422 2544 1480 2550
rect 1422 1856 1480 1862
rect 1422 1822 1434 1856
rect 1422 1816 1480 1822
rect 1830 1514 1888 1520
rect 1830 1480 1842 1514
rect 1830 1474 1888 1480
rect 1398 728 1456 734
rect 1398 694 1410 728
rect 1398 688 1456 694
rect 78 576 136 582
rect 498 576 556 582
rect 78 542 90 576
rect 498 542 510 576
rect 78 536 136 542
rect 498 536 556 542
rect 78 66 136 72
rect 498 66 556 72
rect 78 32 90 66
rect 498 32 510 66
rect 78 26 136 32
rect 498 26 556 32
rect 1398 0 1456 6
rect 1830 4 1888 10
rect 1398 -34 1410 0
rect 1830 -30 1842 4
rect 1398 -40 1456 -34
rect 1830 -36 1888 -30
use sky130_fd_pr__nfet_01v8_ATLS57  XM1
timestamp 1762969946
transform 1 0 107 0 1 304
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_XGSNAL  XM2
timestamp 1762969946
transform 1 0 1451 0 1 2203
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_ATLS57  XM3
timestamp 1762969946
transform 1 0 527 0 1 304
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_XGSNAL  XM4
timestamp 1762969946
transform 1 0 1427 0 1 347
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_KBNS5F  XM5
timestamp 1762969946
transform 1 0 1859 0 1 742
box -211 -910 211 910
<< end >>
